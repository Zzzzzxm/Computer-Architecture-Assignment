
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h19e75bda;
    ram_cell[       1] = 32'h0;  // 32'hbcae6c97;
    ram_cell[       2] = 32'h0;  // 32'he04f1a35;
    ram_cell[       3] = 32'h0;  // 32'h63ef88a9;
    ram_cell[       4] = 32'h0;  // 32'hede79892;
    ram_cell[       5] = 32'h0;  // 32'h5136f6a6;
    ram_cell[       6] = 32'h0;  // 32'hea7ddd4b;
    ram_cell[       7] = 32'h0;  // 32'he7ceb962;
    ram_cell[       8] = 32'h0;  // 32'h1fd332a0;
    ram_cell[       9] = 32'h0;  // 32'h8a93ead2;
    ram_cell[      10] = 32'h0;  // 32'h6911bdf7;
    ram_cell[      11] = 32'h0;  // 32'ha43e04af;
    ram_cell[      12] = 32'h0;  // 32'h8641a381;
    ram_cell[      13] = 32'h0;  // 32'h31677c34;
    ram_cell[      14] = 32'h0;  // 32'hf68da245;
    ram_cell[      15] = 32'h0;  // 32'h9f6049cf;
    ram_cell[      16] = 32'h0;  // 32'h812cccba;
    ram_cell[      17] = 32'h0;  // 32'h1bd64f2b;
    ram_cell[      18] = 32'h0;  // 32'h5c7c8db9;
    ram_cell[      19] = 32'h0;  // 32'hb41f38b3;
    ram_cell[      20] = 32'h0;  // 32'h58676c38;
    ram_cell[      21] = 32'h0;  // 32'h758b8324;
    ram_cell[      22] = 32'h0;  // 32'hd4496bd2;
    ram_cell[      23] = 32'h0;  // 32'h61dd5b3d;
    ram_cell[      24] = 32'h0;  // 32'he44356e5;
    ram_cell[      25] = 32'h0;  // 32'h2a6833b1;
    ram_cell[      26] = 32'h0;  // 32'h572d514b;
    ram_cell[      27] = 32'h0;  // 32'h1710f496;
    ram_cell[      28] = 32'h0;  // 32'h19344585;
    ram_cell[      29] = 32'h0;  // 32'h93abd5f6;
    ram_cell[      30] = 32'h0;  // 32'h0bad06d4;
    ram_cell[      31] = 32'h0;  // 32'hc400258a;
    ram_cell[      32] = 32'h0;  // 32'h3aae5a0a;
    ram_cell[      33] = 32'h0;  // 32'h01401cee;
    ram_cell[      34] = 32'h0;  // 32'hd4d96944;
    ram_cell[      35] = 32'h0;  // 32'hc3a0811c;
    ram_cell[      36] = 32'h0;  // 32'h4c4f6d4c;
    ram_cell[      37] = 32'h0;  // 32'hc267e78d;
    ram_cell[      38] = 32'h0;  // 32'hd88df09e;
    ram_cell[      39] = 32'h0;  // 32'hb9d4c308;
    ram_cell[      40] = 32'h0;  // 32'hf901133a;
    ram_cell[      41] = 32'h0;  // 32'h289aef18;
    ram_cell[      42] = 32'h0;  // 32'h3f322be4;
    ram_cell[      43] = 32'h0;  // 32'h485a00df;
    ram_cell[      44] = 32'h0;  // 32'h9b936730;
    ram_cell[      45] = 32'h0;  // 32'hc5f2bcdc;
    ram_cell[      46] = 32'h0;  // 32'hc91d8d75;
    ram_cell[      47] = 32'h0;  // 32'h0de6dedb;
    ram_cell[      48] = 32'h0;  // 32'h25fe418d;
    ram_cell[      49] = 32'h0;  // 32'h83000bbd;
    ram_cell[      50] = 32'h0;  // 32'h3af70439;
    ram_cell[      51] = 32'h0;  // 32'h97d92712;
    ram_cell[      52] = 32'h0;  // 32'hd98536a4;
    ram_cell[      53] = 32'h0;  // 32'h165b79e7;
    ram_cell[      54] = 32'h0;  // 32'h3e0bb0bd;
    ram_cell[      55] = 32'h0;  // 32'h1bbce1e9;
    ram_cell[      56] = 32'h0;  // 32'h0e524b8f;
    ram_cell[      57] = 32'h0;  // 32'h50b52d23;
    ram_cell[      58] = 32'h0;  // 32'h2a260f5e;
    ram_cell[      59] = 32'h0;  // 32'h9e5ae6e3;
    ram_cell[      60] = 32'h0;  // 32'h2c2c4f46;
    ram_cell[      61] = 32'h0;  // 32'ha98b48ea;
    ram_cell[      62] = 32'h0;  // 32'h88e44e0f;
    ram_cell[      63] = 32'h0;  // 32'h4f42ba10;
    ram_cell[      64] = 32'h0;  // 32'h000cacc8;
    ram_cell[      65] = 32'h0;  // 32'h6f984614;
    ram_cell[      66] = 32'h0;  // 32'hbf0d1d3e;
    ram_cell[      67] = 32'h0;  // 32'h73ea7c75;
    ram_cell[      68] = 32'h0;  // 32'ha1a6489b;
    ram_cell[      69] = 32'h0;  // 32'h65eb1184;
    ram_cell[      70] = 32'h0;  // 32'ha6012070;
    ram_cell[      71] = 32'h0;  // 32'h54648a7b;
    ram_cell[      72] = 32'h0;  // 32'h61f9ec9e;
    ram_cell[      73] = 32'h0;  // 32'h723093e0;
    ram_cell[      74] = 32'h0;  // 32'h9278d0a5;
    ram_cell[      75] = 32'h0;  // 32'h41f70410;
    ram_cell[      76] = 32'h0;  // 32'h784dfd89;
    ram_cell[      77] = 32'h0;  // 32'h2f623773;
    ram_cell[      78] = 32'h0;  // 32'hbb9731ad;
    ram_cell[      79] = 32'h0;  // 32'h624223b8;
    ram_cell[      80] = 32'h0;  // 32'h23f9722c;
    ram_cell[      81] = 32'h0;  // 32'h218d13a5;
    ram_cell[      82] = 32'h0;  // 32'h992c5b2d;
    ram_cell[      83] = 32'h0;  // 32'h983c09c2;
    ram_cell[      84] = 32'h0;  // 32'heffea89d;
    ram_cell[      85] = 32'h0;  // 32'he9a410b0;
    ram_cell[      86] = 32'h0;  // 32'h1d0e930b;
    ram_cell[      87] = 32'h0;  // 32'h4f5cf6ca;
    ram_cell[      88] = 32'h0;  // 32'hb183b825;
    ram_cell[      89] = 32'h0;  // 32'h4cf0d04e;
    ram_cell[      90] = 32'h0;  // 32'hf4bbdee9;
    ram_cell[      91] = 32'h0;  // 32'h6d176b12;
    ram_cell[      92] = 32'h0;  // 32'hddacaa4b;
    ram_cell[      93] = 32'h0;  // 32'h26a4cb90;
    ram_cell[      94] = 32'h0;  // 32'h5e71f680;
    ram_cell[      95] = 32'h0;  // 32'h770ccdf9;
    ram_cell[      96] = 32'h0;  // 32'h0212ec55;
    ram_cell[      97] = 32'h0;  // 32'h76b01fd8;
    ram_cell[      98] = 32'h0;  // 32'hb136c191;
    ram_cell[      99] = 32'h0;  // 32'h8651c7b8;
    ram_cell[     100] = 32'h0;  // 32'he752e96c;
    ram_cell[     101] = 32'h0;  // 32'hdd068e06;
    ram_cell[     102] = 32'h0;  // 32'hc0500cfc;
    ram_cell[     103] = 32'h0;  // 32'h8627c88a;
    ram_cell[     104] = 32'h0;  // 32'h83381a9d;
    ram_cell[     105] = 32'h0;  // 32'heb4538d6;
    ram_cell[     106] = 32'h0;  // 32'h45306ce4;
    ram_cell[     107] = 32'h0;  // 32'h5b3fb660;
    ram_cell[     108] = 32'h0;  // 32'h82d0ff17;
    ram_cell[     109] = 32'h0;  // 32'h156b42eb;
    ram_cell[     110] = 32'h0;  // 32'h5dc84f44;
    ram_cell[     111] = 32'h0;  // 32'h1fba8cbb;
    ram_cell[     112] = 32'h0;  // 32'h8b004e9c;
    ram_cell[     113] = 32'h0;  // 32'hb62c8413;
    ram_cell[     114] = 32'h0;  // 32'h5994a1bc;
    ram_cell[     115] = 32'h0;  // 32'hd0dc7fdc;
    ram_cell[     116] = 32'h0;  // 32'hb5729549;
    ram_cell[     117] = 32'h0;  // 32'h8ecc4cdd;
    ram_cell[     118] = 32'h0;  // 32'hb665c409;
    ram_cell[     119] = 32'h0;  // 32'hc74de3fc;
    ram_cell[     120] = 32'h0;  // 32'h20851d83;
    ram_cell[     121] = 32'h0;  // 32'h15f627db;
    ram_cell[     122] = 32'h0;  // 32'ha63eb7e1;
    ram_cell[     123] = 32'h0;  // 32'hd86da82b;
    ram_cell[     124] = 32'h0;  // 32'h86a97269;
    ram_cell[     125] = 32'h0;  // 32'h6c10021f;
    ram_cell[     126] = 32'h0;  // 32'hcddad150;
    ram_cell[     127] = 32'h0;  // 32'h99368dc2;
    ram_cell[     128] = 32'h0;  // 32'h0dac4eba;
    ram_cell[     129] = 32'h0;  // 32'h31159370;
    ram_cell[     130] = 32'h0;  // 32'h66e064e2;
    ram_cell[     131] = 32'h0;  // 32'h976abcdb;
    ram_cell[     132] = 32'h0;  // 32'h9f0bf972;
    ram_cell[     133] = 32'h0;  // 32'hbfabbc60;
    ram_cell[     134] = 32'h0;  // 32'h3378c599;
    ram_cell[     135] = 32'h0;  // 32'he8dd4146;
    ram_cell[     136] = 32'h0;  // 32'h5dae57b9;
    ram_cell[     137] = 32'h0;  // 32'h432e7742;
    ram_cell[     138] = 32'h0;  // 32'h3d5942f3;
    ram_cell[     139] = 32'h0;  // 32'h29480f95;
    ram_cell[     140] = 32'h0;  // 32'h96de1ccc;
    ram_cell[     141] = 32'h0;  // 32'h28b1e4e1;
    ram_cell[     142] = 32'h0;  // 32'h1fedd69a;
    ram_cell[     143] = 32'h0;  // 32'hbf8f0552;
    ram_cell[     144] = 32'h0;  // 32'h862e9e70;
    ram_cell[     145] = 32'h0;  // 32'hb71e75fe;
    ram_cell[     146] = 32'h0;  // 32'he424e9eb;
    ram_cell[     147] = 32'h0;  // 32'hbf5c3620;
    ram_cell[     148] = 32'h0;  // 32'h7e79b10e;
    ram_cell[     149] = 32'h0;  // 32'h4f1b29b2;
    ram_cell[     150] = 32'h0;  // 32'h28f1e837;
    ram_cell[     151] = 32'h0;  // 32'he3197426;
    ram_cell[     152] = 32'h0;  // 32'h0dff53bf;
    ram_cell[     153] = 32'h0;  // 32'h357605f2;
    ram_cell[     154] = 32'h0;  // 32'h2306eb98;
    ram_cell[     155] = 32'h0;  // 32'h3e01951c;
    ram_cell[     156] = 32'h0;  // 32'h963c9b3a;
    ram_cell[     157] = 32'h0;  // 32'h01cb0a6f;
    ram_cell[     158] = 32'h0;  // 32'ha8489d5d;
    ram_cell[     159] = 32'h0;  // 32'h4a45e978;
    ram_cell[     160] = 32'h0;  // 32'hc84145d5;
    ram_cell[     161] = 32'h0;  // 32'h790bbbaa;
    ram_cell[     162] = 32'h0;  // 32'hf7ca13b1;
    ram_cell[     163] = 32'h0;  // 32'h7db7a3ee;
    ram_cell[     164] = 32'h0;  // 32'hf2157ce8;
    ram_cell[     165] = 32'h0;  // 32'h93765257;
    ram_cell[     166] = 32'h0;  // 32'ha811f859;
    ram_cell[     167] = 32'h0;  // 32'h90b56be8;
    ram_cell[     168] = 32'h0;  // 32'h021e7e5d;
    ram_cell[     169] = 32'h0;  // 32'hfff4775a;
    ram_cell[     170] = 32'h0;  // 32'h40a9b604;
    ram_cell[     171] = 32'h0;  // 32'h7050a2b1;
    ram_cell[     172] = 32'h0;  // 32'h58ef2b95;
    ram_cell[     173] = 32'h0;  // 32'h3614ef79;
    ram_cell[     174] = 32'h0;  // 32'h324b4ac7;
    ram_cell[     175] = 32'h0;  // 32'hefb31381;
    ram_cell[     176] = 32'h0;  // 32'h57d77366;
    ram_cell[     177] = 32'h0;  // 32'heacdc5f3;
    ram_cell[     178] = 32'h0;  // 32'h753d6e2a;
    ram_cell[     179] = 32'h0;  // 32'hdc62ab1d;
    ram_cell[     180] = 32'h0;  // 32'hd54129af;
    ram_cell[     181] = 32'h0;  // 32'h9484b490;
    ram_cell[     182] = 32'h0;  // 32'h34e214d8;
    ram_cell[     183] = 32'h0;  // 32'h7c56c81e;
    ram_cell[     184] = 32'h0;  // 32'h8986513a;
    ram_cell[     185] = 32'h0;  // 32'h4a13e690;
    ram_cell[     186] = 32'h0;  // 32'hb10b1bf1;
    ram_cell[     187] = 32'h0;  // 32'h3af8c1ef;
    ram_cell[     188] = 32'h0;  // 32'h3f5b7ada;
    ram_cell[     189] = 32'h0;  // 32'ha1b953fd;
    ram_cell[     190] = 32'h0;  // 32'h80f414d0;
    ram_cell[     191] = 32'h0;  // 32'h6b5d12ef;
    ram_cell[     192] = 32'h0;  // 32'h560333bf;
    ram_cell[     193] = 32'h0;  // 32'h9e01c771;
    ram_cell[     194] = 32'h0;  // 32'he19fd3dd;
    ram_cell[     195] = 32'h0;  // 32'h4af85379;
    ram_cell[     196] = 32'h0;  // 32'hb186cdca;
    ram_cell[     197] = 32'h0;  // 32'h2ca9ef9c;
    ram_cell[     198] = 32'h0;  // 32'hae27748a;
    ram_cell[     199] = 32'h0;  // 32'hc566aa7b;
    ram_cell[     200] = 32'h0;  // 32'hc04f4bcc;
    ram_cell[     201] = 32'h0;  // 32'hdca2fe1d;
    ram_cell[     202] = 32'h0;  // 32'hfc916b44;
    ram_cell[     203] = 32'h0;  // 32'hdd966dc9;
    ram_cell[     204] = 32'h0;  // 32'h626e10d2;
    ram_cell[     205] = 32'h0;  // 32'he483e48f;
    ram_cell[     206] = 32'h0;  // 32'hf510dc46;
    ram_cell[     207] = 32'h0;  // 32'h312a0570;
    ram_cell[     208] = 32'h0;  // 32'ha1832de8;
    ram_cell[     209] = 32'h0;  // 32'hc7c7abda;
    ram_cell[     210] = 32'h0;  // 32'hbbb61505;
    ram_cell[     211] = 32'h0;  // 32'hd808a9d5;
    ram_cell[     212] = 32'h0;  // 32'h6776496c;
    ram_cell[     213] = 32'h0;  // 32'h141c7967;
    ram_cell[     214] = 32'h0;  // 32'h664ee416;
    ram_cell[     215] = 32'h0;  // 32'h19291357;
    ram_cell[     216] = 32'h0;  // 32'h1fa82f1b;
    ram_cell[     217] = 32'h0;  // 32'hf22cac8b;
    ram_cell[     218] = 32'h0;  // 32'hd1b09633;
    ram_cell[     219] = 32'h0;  // 32'h51b5c7c9;
    ram_cell[     220] = 32'h0;  // 32'h5ed8ffac;
    ram_cell[     221] = 32'h0;  // 32'h729f1ba9;
    ram_cell[     222] = 32'h0;  // 32'h7dfb1f87;
    ram_cell[     223] = 32'h0;  // 32'h95c56ec7;
    ram_cell[     224] = 32'h0;  // 32'hb6da90e3;
    ram_cell[     225] = 32'h0;  // 32'h4360114e;
    ram_cell[     226] = 32'h0;  // 32'h01307aac;
    ram_cell[     227] = 32'h0;  // 32'h1b660c30;
    ram_cell[     228] = 32'h0;  // 32'h7224306a;
    ram_cell[     229] = 32'h0;  // 32'hd77114ee;
    ram_cell[     230] = 32'h0;  // 32'h2f6f4893;
    ram_cell[     231] = 32'h0;  // 32'h0616de09;
    ram_cell[     232] = 32'h0;  // 32'he6be07a6;
    ram_cell[     233] = 32'h0;  // 32'h83d473a4;
    ram_cell[     234] = 32'h0;  // 32'hf0a594c3;
    ram_cell[     235] = 32'h0;  // 32'h6ca60291;
    ram_cell[     236] = 32'h0;  // 32'h075cf3bb;
    ram_cell[     237] = 32'h0;  // 32'h580d1748;
    ram_cell[     238] = 32'h0;  // 32'hef3814e4;
    ram_cell[     239] = 32'h0;  // 32'ha8fce302;
    ram_cell[     240] = 32'h0;  // 32'h1af0e321;
    ram_cell[     241] = 32'h0;  // 32'hbbd63c43;
    ram_cell[     242] = 32'h0;  // 32'h2c48ba60;
    ram_cell[     243] = 32'h0;  // 32'h238312d3;
    ram_cell[     244] = 32'h0;  // 32'h894ebb5d;
    ram_cell[     245] = 32'h0;  // 32'h31024ebd;
    ram_cell[     246] = 32'h0;  // 32'hebbc05d0;
    ram_cell[     247] = 32'h0;  // 32'h95bfed81;
    ram_cell[     248] = 32'h0;  // 32'h99f05bc2;
    ram_cell[     249] = 32'h0;  // 32'hc756007c;
    ram_cell[     250] = 32'h0;  // 32'hcf932854;
    ram_cell[     251] = 32'h0;  // 32'h34b4e99a;
    ram_cell[     252] = 32'h0;  // 32'ha4850568;
    ram_cell[     253] = 32'h0;  // 32'h89c3e879;
    ram_cell[     254] = 32'h0;  // 32'h31c4a14b;
    ram_cell[     255] = 32'h0;  // 32'h01e9f766;
    // src matrix A
    ram_cell[     256] = 32'h8cb009aa;
    ram_cell[     257] = 32'hae000e9e;
    ram_cell[     258] = 32'h7d23a9d3;
    ram_cell[     259] = 32'h95522eee;
    ram_cell[     260] = 32'h2bb6fa2c;
    ram_cell[     261] = 32'he0fd09f9;
    ram_cell[     262] = 32'h49c2037a;
    ram_cell[     263] = 32'h9360db3e;
    ram_cell[     264] = 32'h53b6adb2;
    ram_cell[     265] = 32'h05139a49;
    ram_cell[     266] = 32'hada10c92;
    ram_cell[     267] = 32'hbce36f7a;
    ram_cell[     268] = 32'h574f28d4;
    ram_cell[     269] = 32'h23acb659;
    ram_cell[     270] = 32'he9952eaa;
    ram_cell[     271] = 32'hc9ba89f4;
    ram_cell[     272] = 32'h7e39a13e;
    ram_cell[     273] = 32'h2a4fb2cd;
    ram_cell[     274] = 32'hb837e25e;
    ram_cell[     275] = 32'ha0405d29;
    ram_cell[     276] = 32'hab46f683;
    ram_cell[     277] = 32'h768c4b8a;
    ram_cell[     278] = 32'h51eef38b;
    ram_cell[     279] = 32'h1ae648d5;
    ram_cell[     280] = 32'h1d4932dd;
    ram_cell[     281] = 32'h146b24d8;
    ram_cell[     282] = 32'he1ff589e;
    ram_cell[     283] = 32'h52479983;
    ram_cell[     284] = 32'h465b6dfe;
    ram_cell[     285] = 32'hfcfc4805;
    ram_cell[     286] = 32'h4452f4a6;
    ram_cell[     287] = 32'h12538653;
    ram_cell[     288] = 32'h43f0cef8;
    ram_cell[     289] = 32'h6c033757;
    ram_cell[     290] = 32'h43f01772;
    ram_cell[     291] = 32'hcb717713;
    ram_cell[     292] = 32'h4a550981;
    ram_cell[     293] = 32'h203e7643;
    ram_cell[     294] = 32'h57f10eab;
    ram_cell[     295] = 32'hb4490864;
    ram_cell[     296] = 32'hc1c54fa4;
    ram_cell[     297] = 32'h0b0954ac;
    ram_cell[     298] = 32'h6b24e0a0;
    ram_cell[     299] = 32'h69291b77;
    ram_cell[     300] = 32'ha26cc6c9;
    ram_cell[     301] = 32'hf4a6f0ff;
    ram_cell[     302] = 32'h516b97e1;
    ram_cell[     303] = 32'hf904c51d;
    ram_cell[     304] = 32'h15ba6e13;
    ram_cell[     305] = 32'hec1fad46;
    ram_cell[     306] = 32'h3cad1a25;
    ram_cell[     307] = 32'h4a8eff31;
    ram_cell[     308] = 32'h8d452c71;
    ram_cell[     309] = 32'hfdc1046d;
    ram_cell[     310] = 32'hda10f2b7;
    ram_cell[     311] = 32'h5d8f4817;
    ram_cell[     312] = 32'h9da21617;
    ram_cell[     313] = 32'h7373a0b1;
    ram_cell[     314] = 32'h0eb7da31;
    ram_cell[     315] = 32'h0ac3876d;
    ram_cell[     316] = 32'h0158074c;
    ram_cell[     317] = 32'h664e3778;
    ram_cell[     318] = 32'ha78650be;
    ram_cell[     319] = 32'h8eaa96ce;
    ram_cell[     320] = 32'he0801515;
    ram_cell[     321] = 32'h54d76e60;
    ram_cell[     322] = 32'ha9c1604f;
    ram_cell[     323] = 32'h2d3f7da3;
    ram_cell[     324] = 32'h13bfa08c;
    ram_cell[     325] = 32'h88561421;
    ram_cell[     326] = 32'h89c64e31;
    ram_cell[     327] = 32'h6dc07816;
    ram_cell[     328] = 32'h6717031e;
    ram_cell[     329] = 32'h1f27c9d3;
    ram_cell[     330] = 32'h18bd3bf1;
    ram_cell[     331] = 32'h3dba6ec2;
    ram_cell[     332] = 32'h7c994cbc;
    ram_cell[     333] = 32'hf7a7affb;
    ram_cell[     334] = 32'h17355ae5;
    ram_cell[     335] = 32'hccd25e80;
    ram_cell[     336] = 32'he8b2644a;
    ram_cell[     337] = 32'hc744ecf4;
    ram_cell[     338] = 32'h1039d783;
    ram_cell[     339] = 32'h43da5f89;
    ram_cell[     340] = 32'hd03a62f6;
    ram_cell[     341] = 32'hd262f64f;
    ram_cell[     342] = 32'h552e20bd;
    ram_cell[     343] = 32'h2284202e;
    ram_cell[     344] = 32'h0ca210d1;
    ram_cell[     345] = 32'h35393961;
    ram_cell[     346] = 32'h492b97fa;
    ram_cell[     347] = 32'h16452d36;
    ram_cell[     348] = 32'had456c5a;
    ram_cell[     349] = 32'hd9507025;
    ram_cell[     350] = 32'h38a98ee3;
    ram_cell[     351] = 32'ha2faa068;
    ram_cell[     352] = 32'h8d5d5b30;
    ram_cell[     353] = 32'hb196792e;
    ram_cell[     354] = 32'h709e14f5;
    ram_cell[     355] = 32'h9bce1937;
    ram_cell[     356] = 32'h3699602f;
    ram_cell[     357] = 32'h1a0b29ac;
    ram_cell[     358] = 32'he90fca74;
    ram_cell[     359] = 32'h1e9c28e4;
    ram_cell[     360] = 32'hfcff3bfa;
    ram_cell[     361] = 32'ha7e34833;
    ram_cell[     362] = 32'h740961be;
    ram_cell[     363] = 32'h1b67cdd3;
    ram_cell[     364] = 32'h84e6e663;
    ram_cell[     365] = 32'h622e45e9;
    ram_cell[     366] = 32'h04598918;
    ram_cell[     367] = 32'h8e1bb18f;
    ram_cell[     368] = 32'hde14e757;
    ram_cell[     369] = 32'hba6fd7e7;
    ram_cell[     370] = 32'h548be715;
    ram_cell[     371] = 32'h30a626d0;
    ram_cell[     372] = 32'h753e09df;
    ram_cell[     373] = 32'h7d1707cc;
    ram_cell[     374] = 32'h0f8bb8db;
    ram_cell[     375] = 32'hf00ef28a;
    ram_cell[     376] = 32'h6e18819a;
    ram_cell[     377] = 32'h5ceb7325;
    ram_cell[     378] = 32'h2196d481;
    ram_cell[     379] = 32'h85978b2a;
    ram_cell[     380] = 32'he731f097;
    ram_cell[     381] = 32'h5a94ae27;
    ram_cell[     382] = 32'h9f5bf5b2;
    ram_cell[     383] = 32'h9eeadb07;
    ram_cell[     384] = 32'h6cdc150b;
    ram_cell[     385] = 32'hd3a8363f;
    ram_cell[     386] = 32'haa7cf09e;
    ram_cell[     387] = 32'hf047c278;
    ram_cell[     388] = 32'ha21ab4cd;
    ram_cell[     389] = 32'hc579d3d4;
    ram_cell[     390] = 32'ha3a8e316;
    ram_cell[     391] = 32'h1970169d;
    ram_cell[     392] = 32'hb0ea80c0;
    ram_cell[     393] = 32'haf27be0f;
    ram_cell[     394] = 32'h88724ad3;
    ram_cell[     395] = 32'h97a17f65;
    ram_cell[     396] = 32'hd5189af4;
    ram_cell[     397] = 32'h17959bcc;
    ram_cell[     398] = 32'h96178b82;
    ram_cell[     399] = 32'h34e3a1b7;
    ram_cell[     400] = 32'h60892130;
    ram_cell[     401] = 32'h18821109;
    ram_cell[     402] = 32'hf9bff4a3;
    ram_cell[     403] = 32'h1718d8a5;
    ram_cell[     404] = 32'h36c9459b;
    ram_cell[     405] = 32'h5401752c;
    ram_cell[     406] = 32'hdde0d27f;
    ram_cell[     407] = 32'h71ff6f15;
    ram_cell[     408] = 32'h6e1b46a3;
    ram_cell[     409] = 32'h94ec1465;
    ram_cell[     410] = 32'h78a38950;
    ram_cell[     411] = 32'h16ca58ed;
    ram_cell[     412] = 32'h6b3f3dec;
    ram_cell[     413] = 32'h076f16c7;
    ram_cell[     414] = 32'he59bd356;
    ram_cell[     415] = 32'hdc4e7d3a;
    ram_cell[     416] = 32'h573537df;
    ram_cell[     417] = 32'h325f9df9;
    ram_cell[     418] = 32'hc99a1cfc;
    ram_cell[     419] = 32'hdb1abf4d;
    ram_cell[     420] = 32'h1274cd67;
    ram_cell[     421] = 32'hb0e7ff0e;
    ram_cell[     422] = 32'hb149cd2d;
    ram_cell[     423] = 32'ha6c39e4d;
    ram_cell[     424] = 32'h9349eb14;
    ram_cell[     425] = 32'h2f2a7cf0;
    ram_cell[     426] = 32'h604b0004;
    ram_cell[     427] = 32'h1fa264ec;
    ram_cell[     428] = 32'h3575bb18;
    ram_cell[     429] = 32'h5df8ecc0;
    ram_cell[     430] = 32'hd1922458;
    ram_cell[     431] = 32'hd80911a8;
    ram_cell[     432] = 32'h6f859839;
    ram_cell[     433] = 32'hf07f8da1;
    ram_cell[     434] = 32'h240e54ac;
    ram_cell[     435] = 32'hce8f4f5b;
    ram_cell[     436] = 32'h10e639c3;
    ram_cell[     437] = 32'h91b36930;
    ram_cell[     438] = 32'ha5e24fe0;
    ram_cell[     439] = 32'hd31b17a3;
    ram_cell[     440] = 32'h55c779ce;
    ram_cell[     441] = 32'h60e7e099;
    ram_cell[     442] = 32'hb3ce62f1;
    ram_cell[     443] = 32'hcac834cf;
    ram_cell[     444] = 32'h5aa79b77;
    ram_cell[     445] = 32'hd2cda3c2;
    ram_cell[     446] = 32'h02dc29d8;
    ram_cell[     447] = 32'he2f15345;
    ram_cell[     448] = 32'h7e4fbb72;
    ram_cell[     449] = 32'he528a20a;
    ram_cell[     450] = 32'h9219fec3;
    ram_cell[     451] = 32'h7772d0ed;
    ram_cell[     452] = 32'hfc862fb0;
    ram_cell[     453] = 32'h0f2ef809;
    ram_cell[     454] = 32'h29d945f0;
    ram_cell[     455] = 32'h14867ff1;
    ram_cell[     456] = 32'hbbe581d9;
    ram_cell[     457] = 32'haeb35d4b;
    ram_cell[     458] = 32'h04b585ff;
    ram_cell[     459] = 32'hc312ac24;
    ram_cell[     460] = 32'hf73f00ed;
    ram_cell[     461] = 32'he494db7b;
    ram_cell[     462] = 32'h7f79a68b;
    ram_cell[     463] = 32'hccdc44e6;
    ram_cell[     464] = 32'hcbcc346b;
    ram_cell[     465] = 32'hc24b18a2;
    ram_cell[     466] = 32'h7f7238c7;
    ram_cell[     467] = 32'hbbd9cbd3;
    ram_cell[     468] = 32'h166836c6;
    ram_cell[     469] = 32'ha3ce5985;
    ram_cell[     470] = 32'hd9c8cd08;
    ram_cell[     471] = 32'haf9cd0e4;
    ram_cell[     472] = 32'h7dbdc5f0;
    ram_cell[     473] = 32'h6fbe31a7;
    ram_cell[     474] = 32'h6f79884c;
    ram_cell[     475] = 32'hfb66d442;
    ram_cell[     476] = 32'h7f3c27d2;
    ram_cell[     477] = 32'hb3a3007e;
    ram_cell[     478] = 32'h69884d1d;
    ram_cell[     479] = 32'hb6c1c89e;
    ram_cell[     480] = 32'h180ccea6;
    ram_cell[     481] = 32'h17408741;
    ram_cell[     482] = 32'h0530c8f4;
    ram_cell[     483] = 32'h3270e2cf;
    ram_cell[     484] = 32'h370fcd5b;
    ram_cell[     485] = 32'h94943f92;
    ram_cell[     486] = 32'h09a17bf1;
    ram_cell[     487] = 32'h786d96c3;
    ram_cell[     488] = 32'he5e67ace;
    ram_cell[     489] = 32'h56b90af0;
    ram_cell[     490] = 32'he5224529;
    ram_cell[     491] = 32'h886d2c7c;
    ram_cell[     492] = 32'hbf82657f;
    ram_cell[     493] = 32'hb6437c56;
    ram_cell[     494] = 32'h9087b1aa;
    ram_cell[     495] = 32'h6400bd5e;
    ram_cell[     496] = 32'h101d3b5c;
    ram_cell[     497] = 32'h08bfbbbd;
    ram_cell[     498] = 32'h2a5228c5;
    ram_cell[     499] = 32'hb81a89cd;
    ram_cell[     500] = 32'h54b3329e;
    ram_cell[     501] = 32'h31fddfbb;
    ram_cell[     502] = 32'h6c9ab717;
    ram_cell[     503] = 32'he0b4b552;
    ram_cell[     504] = 32'h02c61500;
    ram_cell[     505] = 32'h24f0feb5;
    ram_cell[     506] = 32'h7adb7fdf;
    ram_cell[     507] = 32'hcdba3ab0;
    ram_cell[     508] = 32'hd1158b9e;
    ram_cell[     509] = 32'hb2e8e55f;
    ram_cell[     510] = 32'h37eca776;
    ram_cell[     511] = 32'h05092089;
    // src matrix B
    ram_cell[     512] = 32'h301b88c6;
    ram_cell[     513] = 32'hb8fc5ce1;
    ram_cell[     514] = 32'he5d86975;
    ram_cell[     515] = 32'hc4d42834;
    ram_cell[     516] = 32'h4cfed510;
    ram_cell[     517] = 32'he4b6f8b4;
    ram_cell[     518] = 32'hd1400607;
    ram_cell[     519] = 32'hf90dc96b;
    ram_cell[     520] = 32'h20dde628;
    ram_cell[     521] = 32'h2c711f74;
    ram_cell[     522] = 32'hc41a503c;
    ram_cell[     523] = 32'h1d3ccfb4;
    ram_cell[     524] = 32'h55145ac9;
    ram_cell[     525] = 32'hac7050b9;
    ram_cell[     526] = 32'hb221d1c3;
    ram_cell[     527] = 32'h41676d27;
    ram_cell[     528] = 32'ha6706eb9;
    ram_cell[     529] = 32'h91e9fd73;
    ram_cell[     530] = 32'hc7dc74d0;
    ram_cell[     531] = 32'h756de3d9;
    ram_cell[     532] = 32'h5b7ac7f3;
    ram_cell[     533] = 32'hd3494006;
    ram_cell[     534] = 32'hdb4519d7;
    ram_cell[     535] = 32'h32d42c38;
    ram_cell[     536] = 32'h829d9336;
    ram_cell[     537] = 32'h23a12e8b;
    ram_cell[     538] = 32'he76677cc;
    ram_cell[     539] = 32'h449551f9;
    ram_cell[     540] = 32'hdf34316e;
    ram_cell[     541] = 32'h37b8837f;
    ram_cell[     542] = 32'h1fe11c06;
    ram_cell[     543] = 32'he78c9c6d;
    ram_cell[     544] = 32'h58f70e41;
    ram_cell[     545] = 32'h45d7440a;
    ram_cell[     546] = 32'hda8fb88d;
    ram_cell[     547] = 32'h4fb3c199;
    ram_cell[     548] = 32'h7fd9f5e0;
    ram_cell[     549] = 32'hf8cef8be;
    ram_cell[     550] = 32'ha6ab89d2;
    ram_cell[     551] = 32'hc4b9f566;
    ram_cell[     552] = 32'h4214c0d4;
    ram_cell[     553] = 32'h7a063927;
    ram_cell[     554] = 32'h2244d341;
    ram_cell[     555] = 32'h23eb820c;
    ram_cell[     556] = 32'h8297b1a5;
    ram_cell[     557] = 32'hdf833c67;
    ram_cell[     558] = 32'h7907ba1b;
    ram_cell[     559] = 32'ha0ad4f80;
    ram_cell[     560] = 32'hb752bd9d;
    ram_cell[     561] = 32'h7dc245fa;
    ram_cell[     562] = 32'h43ad9f80;
    ram_cell[     563] = 32'h03cff164;
    ram_cell[     564] = 32'ha41a9db4;
    ram_cell[     565] = 32'h7db78b72;
    ram_cell[     566] = 32'h6435d7f1;
    ram_cell[     567] = 32'h5ecb42a2;
    ram_cell[     568] = 32'h8ddb3ce8;
    ram_cell[     569] = 32'h801e483d;
    ram_cell[     570] = 32'h08281ff8;
    ram_cell[     571] = 32'h8d21d5e1;
    ram_cell[     572] = 32'h1c78527d;
    ram_cell[     573] = 32'h27ad5414;
    ram_cell[     574] = 32'h3c405f3c;
    ram_cell[     575] = 32'h32cd9945;
    ram_cell[     576] = 32'hd3097c28;
    ram_cell[     577] = 32'hdd9e4fa3;
    ram_cell[     578] = 32'h1197bf52;
    ram_cell[     579] = 32'h4514c5cc;
    ram_cell[     580] = 32'h73e26906;
    ram_cell[     581] = 32'h5e82e460;
    ram_cell[     582] = 32'hb4bedc3e;
    ram_cell[     583] = 32'hdce04754;
    ram_cell[     584] = 32'hf68fb8e3;
    ram_cell[     585] = 32'h88e0ff1f;
    ram_cell[     586] = 32'hc58f9ff8;
    ram_cell[     587] = 32'h129abb60;
    ram_cell[     588] = 32'h9424c8d9;
    ram_cell[     589] = 32'h71e9fde2;
    ram_cell[     590] = 32'h58a2e6c2;
    ram_cell[     591] = 32'h9c4c79f9;
    ram_cell[     592] = 32'h7ebe3bc9;
    ram_cell[     593] = 32'h9514f735;
    ram_cell[     594] = 32'h3f9532f5;
    ram_cell[     595] = 32'h4c2a6fd5;
    ram_cell[     596] = 32'h3cf30319;
    ram_cell[     597] = 32'hc65344fa;
    ram_cell[     598] = 32'h3c2df191;
    ram_cell[     599] = 32'h4f0346a4;
    ram_cell[     600] = 32'h7f4842ff;
    ram_cell[     601] = 32'h1b9240e4;
    ram_cell[     602] = 32'ha8682f6f;
    ram_cell[     603] = 32'hbb162d3f;
    ram_cell[     604] = 32'h145950f9;
    ram_cell[     605] = 32'h7791af39;
    ram_cell[     606] = 32'h07dd21f4;
    ram_cell[     607] = 32'h882bd657;
    ram_cell[     608] = 32'h3e1fbb99;
    ram_cell[     609] = 32'h11de6da6;
    ram_cell[     610] = 32'h247a1c61;
    ram_cell[     611] = 32'hedfa7f78;
    ram_cell[     612] = 32'h3279e875;
    ram_cell[     613] = 32'h1cbab5c8;
    ram_cell[     614] = 32'h46fec00d;
    ram_cell[     615] = 32'ha18b9c9e;
    ram_cell[     616] = 32'hc621575e;
    ram_cell[     617] = 32'h9e2fd219;
    ram_cell[     618] = 32'hcead5ed9;
    ram_cell[     619] = 32'h51e025e6;
    ram_cell[     620] = 32'h840eb079;
    ram_cell[     621] = 32'h7fa98de0;
    ram_cell[     622] = 32'hd8ced651;
    ram_cell[     623] = 32'hf20b1a08;
    ram_cell[     624] = 32'h318a8e18;
    ram_cell[     625] = 32'h53597f9b;
    ram_cell[     626] = 32'hd5fcaf95;
    ram_cell[     627] = 32'he681eaf5;
    ram_cell[     628] = 32'h3d9bc302;
    ram_cell[     629] = 32'hfffce8ff;
    ram_cell[     630] = 32'heabc471d;
    ram_cell[     631] = 32'h5c357c79;
    ram_cell[     632] = 32'hb180e3c6;
    ram_cell[     633] = 32'h3cd4a558;
    ram_cell[     634] = 32'h02d2980d;
    ram_cell[     635] = 32'h5fe002ed;
    ram_cell[     636] = 32'h06744ff1;
    ram_cell[     637] = 32'h5ff3f26b;
    ram_cell[     638] = 32'h089300c3;
    ram_cell[     639] = 32'h37455195;
    ram_cell[     640] = 32'h37a73875;
    ram_cell[     641] = 32'h587893b2;
    ram_cell[     642] = 32'hb6c1ae04;
    ram_cell[     643] = 32'h9e44f2bd;
    ram_cell[     644] = 32'h3fc88973;
    ram_cell[     645] = 32'hc028a797;
    ram_cell[     646] = 32'hc96b98a5;
    ram_cell[     647] = 32'hc93270a8;
    ram_cell[     648] = 32'h5dedfa5b;
    ram_cell[     649] = 32'hcd0de403;
    ram_cell[     650] = 32'h9d73cc5b;
    ram_cell[     651] = 32'hc07d860d;
    ram_cell[     652] = 32'h6bba7381;
    ram_cell[     653] = 32'h48949f1e;
    ram_cell[     654] = 32'h9cff28fa;
    ram_cell[     655] = 32'ha17f24fe;
    ram_cell[     656] = 32'hbc31a468;
    ram_cell[     657] = 32'hbde8635a;
    ram_cell[     658] = 32'hd66c5ab1;
    ram_cell[     659] = 32'h82ba4e0b;
    ram_cell[     660] = 32'h784f3cda;
    ram_cell[     661] = 32'h2836a0a6;
    ram_cell[     662] = 32'h748fd384;
    ram_cell[     663] = 32'h88e5126e;
    ram_cell[     664] = 32'h755500d4;
    ram_cell[     665] = 32'h1b19c022;
    ram_cell[     666] = 32'h79273139;
    ram_cell[     667] = 32'hb381426a;
    ram_cell[     668] = 32'h0eaf834d;
    ram_cell[     669] = 32'hf578a078;
    ram_cell[     670] = 32'h42888b19;
    ram_cell[     671] = 32'h5caf315b;
    ram_cell[     672] = 32'hdd7ed50d;
    ram_cell[     673] = 32'hf9dcf32a;
    ram_cell[     674] = 32'h17d10b7c;
    ram_cell[     675] = 32'hdbe88b84;
    ram_cell[     676] = 32'h26e44b37;
    ram_cell[     677] = 32'hdcacf55b;
    ram_cell[     678] = 32'h437d7301;
    ram_cell[     679] = 32'h08b265b8;
    ram_cell[     680] = 32'h8840ac9c;
    ram_cell[     681] = 32'h4e6f8291;
    ram_cell[     682] = 32'h6a448423;
    ram_cell[     683] = 32'hdf775b9b;
    ram_cell[     684] = 32'ha014db66;
    ram_cell[     685] = 32'h156c199a;
    ram_cell[     686] = 32'h9d5d3a0a;
    ram_cell[     687] = 32'hce574e46;
    ram_cell[     688] = 32'h7d750eb1;
    ram_cell[     689] = 32'hfa155e8f;
    ram_cell[     690] = 32'h97ad6797;
    ram_cell[     691] = 32'h7ffb141b;
    ram_cell[     692] = 32'he89fad74;
    ram_cell[     693] = 32'h3f6b83a6;
    ram_cell[     694] = 32'hb8ed30cc;
    ram_cell[     695] = 32'he48a7cf7;
    ram_cell[     696] = 32'h0a706776;
    ram_cell[     697] = 32'hfc89c809;
    ram_cell[     698] = 32'he647e9ff;
    ram_cell[     699] = 32'h7538d74c;
    ram_cell[     700] = 32'ha7ddd76f;
    ram_cell[     701] = 32'h0f3e2258;
    ram_cell[     702] = 32'h22e8fbea;
    ram_cell[     703] = 32'he77ceb48;
    ram_cell[     704] = 32'h1cb6c25f;
    ram_cell[     705] = 32'h69378b91;
    ram_cell[     706] = 32'hed26b34c;
    ram_cell[     707] = 32'he159d4a4;
    ram_cell[     708] = 32'h7facd6c7;
    ram_cell[     709] = 32'h4be97794;
    ram_cell[     710] = 32'h018b3e14;
    ram_cell[     711] = 32'h593c43a4;
    ram_cell[     712] = 32'hf14d3ba7;
    ram_cell[     713] = 32'h92e19f8f;
    ram_cell[     714] = 32'hb1b42a20;
    ram_cell[     715] = 32'he2a51a25;
    ram_cell[     716] = 32'h04c9ed39;
    ram_cell[     717] = 32'hc40ed1fe;
    ram_cell[     718] = 32'he090faf4;
    ram_cell[     719] = 32'hdc8dc394;
    ram_cell[     720] = 32'hdeb7f822;
    ram_cell[     721] = 32'h52dd697e;
    ram_cell[     722] = 32'h81269092;
    ram_cell[     723] = 32'h0f9680e2;
    ram_cell[     724] = 32'hc00df85d;
    ram_cell[     725] = 32'ha0057f0a;
    ram_cell[     726] = 32'h2bbb7e4c;
    ram_cell[     727] = 32'hd4ec1a2e;
    ram_cell[     728] = 32'h92707de7;
    ram_cell[     729] = 32'h73a4c1f1;
    ram_cell[     730] = 32'h1d2d1864;
    ram_cell[     731] = 32'h5502e3a2;
    ram_cell[     732] = 32'h9e60f978;
    ram_cell[     733] = 32'h20fe377a;
    ram_cell[     734] = 32'h2de2e169;
    ram_cell[     735] = 32'h49570fcb;
    ram_cell[     736] = 32'h59fd1d27;
    ram_cell[     737] = 32'h929577be;
    ram_cell[     738] = 32'h9cdd6069;
    ram_cell[     739] = 32'hd3c90b88;
    ram_cell[     740] = 32'h9ce86ce1;
    ram_cell[     741] = 32'h27901499;
    ram_cell[     742] = 32'h18100c0d;
    ram_cell[     743] = 32'h01a3e6a4;
    ram_cell[     744] = 32'h4fdf91b8;
    ram_cell[     745] = 32'hc334acdf;
    ram_cell[     746] = 32'h8230e7ae;
    ram_cell[     747] = 32'h2ab7774f;
    ram_cell[     748] = 32'hc5355f1d;
    ram_cell[     749] = 32'h07229884;
    ram_cell[     750] = 32'h2245495c;
    ram_cell[     751] = 32'hb3733577;
    ram_cell[     752] = 32'hcc6ebfb7;
    ram_cell[     753] = 32'h7076bdd7;
    ram_cell[     754] = 32'h5dca198a;
    ram_cell[     755] = 32'h851325dd;
    ram_cell[     756] = 32'hd051515e;
    ram_cell[     757] = 32'hcaa92c8e;
    ram_cell[     758] = 32'haed8d7df;
    ram_cell[     759] = 32'h6d99b833;
    ram_cell[     760] = 32'h1409eb78;
    ram_cell[     761] = 32'h412f65ee;
    ram_cell[     762] = 32'he198d4a7;
    ram_cell[     763] = 32'h8e173e82;
    ram_cell[     764] = 32'h9d0d6eb3;
    ram_cell[     765] = 32'ha5c1705c;
    ram_cell[     766] = 32'h6aab70fb;
    ram_cell[     767] = 32'hd7b6f40d;
end

endmodule

